`define CFG_SYS_FREQ                   50000000
`define CFG_BAUD_RATE                  9600
`define CFG_SAMPLE                     16
